library verilog;
use verilog.vl_types.all;
entity traditional_multiplier16_tb is
end traditional_multiplier16_tb;
